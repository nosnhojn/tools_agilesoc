module myAxiStreamingCgModule
(
  input clk,
  input rst_n,
