  endgroup

endmodule

