module myAxiStreamingCgModule
(
